`timescale 1ns / 1ps
module clock(input  logic clk,
             output logic clk_en);
 //10^8? 
//logic clk_en;

endmodule
